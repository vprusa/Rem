	
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
USE ieee.math_real.ALL;   -- for UNIFORM, TRUNC functions
USE ieee.numeric_std.ALL; -- for TO_UNSIGNED function

use work.vga_controller_cfg.all;

architecture behav of tlv_pc_ifc is 
  signal vga_mode: std_logic_vector(60 downto 0);
  signal red: std_logic_vector(2 downto 0);
  signal green: std_logic_vector(2 downto 0);
  signal blue: std_logic_vector(2 downto 0);
  signal rgb : std_logic_vector(8 downto 0);
  signal rgbMsg : std_logic_vector(8 downto 0);
  signal rgbLvlMsg : std_logic_vector(8 downto 0);
  signal rgbLvlNmb : std_logic_vector(8 downto 0);
  signal rgbf : std_logic_vector(8 downto 0);

  signal vgaRow: std_logic_vector(11 downto 0);
  signal vgaCol: std_logic_vector(11 downto 0);

  signal en_2Hz,en_4Hz, en_8Hz, en_16Hz, en_1MHz, en_20Hz : std_logic;
  signal random_nmb : std_logic_vector(7 downto 0) := (4 => '1',2 => '1',others => '0');
 
  signal digger_clr : std_logic_vector(0 to 1);
  signal current_nmb_index : integer range 0 to 9 := 0;
  signal rom_col : integer range 0 to 32;
 
  type generated_type is array(9 downto 0) of integer range 0 to 9;
  signal generated_rand : generated_type := (others => (integer(0)));
  
  type t_key is (K0,K1,K2,K3,K4,K5,K6,K7,K8,K9,KA,KB,KC,KD,KHASH,KSTAR,NONE);
  signal key_pressed : t_key := NONE; 
  signal key_read : std_logic := '0';
  signal number_pressed : std_logic_vector (3 downto 0) := "1111";
  type t_key_signal_check is array(2 downto 0) of std_logic_vector (3 downto 0);
  type t_text is (NONE,BEFORE_WRITING_NUMBERS,LEVEL_OK,LEVEL_BAD);
  signal text : t_text := NONE; 

  type t_game_states is (WELCOME_SCREEN,WAITING_SCREEN,GEN_NMB, SHOWING_NUMBERS, WRITING_NUMBERS,LEVEL_END_BAD,LEVEL_END_OK,CONFIG_SPEED);
  signal game_state : t_game_states := WELCOME_SCREEN; 
  
	signal game_speed : std_logic_vector(2 downto 0) := "010";
	signal game_level : integer := 1;

	constant MAX_INDEX : integer := 7;
	constant MIN_INDEX : integer := 1;
 
  type pamet_nmb is array(0 to 16*10) of std_logic_vector(0 to 31);
  type pamet_msg is array(0 to 16*5) of std_logic_vector(0 to 319);-- ? 320 ?
   type pamet_lvl is array(0 to 8) of std_logic_vector(0 to 63);-- ? 160 ?

signal rom_lvl: pamet_lvl := ( 
"0001000000011111101000001001111110010000000000000000000000000000",
"0001000000010000001000001001000000010000000000000000000000000000",
"0001000000010000000100010001000000010000000000000000000000000000",
"0001000000011111000100010001111100010000000000000000000000000000",
"0001000000010000000010100001000000010000000000000000000000000000",
"0001000000010000000010100001000000010000000000000000000000000000",
"0001000000010000000001000001000000010000000000000000000000000000",
"0001111110011111100001000001111110011111100000000000000000000000",
(others => '0'));

signal rom_msg: pamet_msg := (
"00100000100111111001000000001111000011110010000010011111100000000000000000000000000111110001111100011111100011110000111100000000000000000000000000111111100011110000000000001111001111111000011000011111001111111000000000000110000100001001111000000000000111110001111110100000100111111010000010011111000111111001111100000100",
"00100000100100000001000000010000100100001011000110010000000000000000000000000000000100001001000010010000000100001001000010000000000001001000000000000100000100001000000000010000100001000000100100010000100001000000000000001001000110001001000100000000000100001001000000110001100100000011000110010000100100000001000010000100",
"00100100100100000001000000010000000100001010101010010000000000000000000000000000000100001001000010010000000100000001000000000000000001001000000000000100000100001000000000010000000001000001000010010000100001000000000000010000100101001001000010000000000100001001000000101010100100000010101010010000100100000001000010000100",
"00100100100111110001000000010000000100001010101010011111000000000000000000000000000111110001111100011111000011000000110000000000000111111100000000000100000100001000000000001100000001000001000010011111000001000000000000010000100101001001000010000000000111110001111100101010100111110010101010011111000111110001111100000100",
"00100100100100000001000000010000000100001010010010010000000000000001111110000000000100000001001000010000000000110000001100000000000010010000000000000100000100001000000000000011000001000001111110010010000001000000000000011111100100101001000010000000000100100001000000100100100100000010010010010000100100000001001000000100",
"00100100100100000001000000010000000100001010010010010000000000000000000000000000000100000001000100010000000000001000000010000000001111111000000000000100000100001000000000000000100001000001000010010001000001000000000000010000100100101001000010000000000100010001000000100100100100000010010010010000100100000001000100000100",
"00101010100100000001000000010000100100001010000010010000000000000000000000000000000100000001000010010000000100001001000010000000000100100000000000000100000100001000000000010000100001000001000010010000100001000000000000010000100100011001000100000000000100001001000000100000100100000010000010010000100100000001000010000100",
"00010001000111111001111110001111000011110010000010011111100000000000000000000000000100000001000010011111100011110000111100000000000100100000000000000100000011110000000000001111000001000001000010010000100001000000000000010000100100001001111000000000000100001001111110100000100111111010000010011111000111111001000010000100",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
"00100000100011110001000010000000001000001000111100010000100000000000000000000000000111110001111100011111100011110000111100000000000000000000000000011111100011110001111100000000000100001001111110010000101111111000000000011111000011110001000010010000100111100000000000000000000000000000000000000000000000000000000000000000",
"00100000100100001001000010000000001000001001000010011000100000000000000000000000000100001001000010010000000100001001000010000000010000010000000000010000000100001001000010000000000110001001000000010000100001000000000000010000100100001001000010011000100100010000000000000000000000000000000000000000000000000000000000000000",
"00010001000100001001000010000000001001001001000010010100100000000000000000000000000100001001000010010000000100000001000000000000001000100000000000010000000100001001000010000000000101001001000000001001000001000000000000010000100100001001000010010100100100001000000000000000000000000000000000000000000000000000000000000000",
"00001010000100001001000010000000001001001001000010010100100000000000000000000000000111110001111100011111000011000000110000000000000101000000000000011111000100001001111100000000000101001001111100000110000001000000000000011111000100001001000010010100100100001000000000000000000000000000000000000000000000000000000000000000",
"00000100000100001001000010000000001001001001000010010010100000000001111110000000000100000001001000010000000000110000001100000000111111111000000000010000000100001001001000000000000100101001000000000110000001000000000000010010000100001001000010010010100100001000000000000000000000000000000000000000000000000000000000000000",
"00000100000100001001000010000000001001001001000010010010100000000000000000000000000100000001000100010000000000001000000010000000000101000000000000010000000100001001000100000000000100101001000000001001000001000000000000010001000100001001000010010010100100001000000000000000000000000000000000000000000000000000000000000000",
"00000100000100001001000010000000001010101001000010010001100000000000000000000000000100000001000010010000000100001001000010000000001000100000000000010000000100001001000010000000000100011001000000010000100001000000000000010000100100001001000010010001100100010000000000000000000000000000000000000000000000000000000000000000",
"00000100000011110000111100000000000100010000111100010000100000000000000000000000000100000001000010011111100011110000111100000000010000010000000000010000000011110001000010000000000100001001111110010000100001000000000000010000100011110000111100010000100111100000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
"00100000100011110001000010000000000100000000111100001111001111111000000000000000000000000001111100011111000111111000111100001111000000000000000000000000001111111000111100000000000011110000111100010000101111111001111100010000100100001001111110000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00100000100100001001000010000000000100000001000010010000100001000000000000000000000000000001000010010000100100000001000010010000100000000010001000000000000001000001000010000000000100001001000010011000100001000000010000011000100100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00001010000100001001000010000000000100000001000010001100000001000000000000000000000000000001111100011111000111110000110000001100000000000001010000000000000001000001000010000000000100000001000010010100100001000000010000010100100100001001111100000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000100000100001001000010000000000100000001000010000011000001000000000000011111100000000001000000010010000100000000001100000011000000001111111110000000000001000001000010000000000100000001000010010010100001000000010000010010100100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000100000100001001000010000000000100000001000010000000100001000000000000000000000000000001000000010001000100000000000010000000100000000001010000000000000001000001000010000000000100000001000010010010100001000000010000010010100100001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000100000011110000111100000000000111111000111100001111000001000000000000000000000000000001000000010000100111111000111100001111000000000010001000000000000001000000111100000000000011110000111100010000100001000001111100010000100011110001111110000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
"00011111000111110001111110001111000011110000000000010000100100001010000010011111000111111001111100001111000000000001111100010000100000000000111100011111000111100001111110011111000000000010000010001111000100001000000000011111000111111010000010011111101000001001111100011111100111110000000000000000000000000000000000000000",
"00010000100100001001000000010000100100001000000000011000100100001011000110010000100100000001000010010000100000000000010000011000100000000001000010010000100100010001000000010000100000000010000010010000100100001000000000010000100100000011000110010000001100011001000010010000000100001000000000000000000000000000000000000000",
"00010000100100001001000000010000000100000000000000010100100100001010101010010000100100000001000010010000000000000000010000010100100000000001000010010000100100001001000000010000100000000001000100010000100100001000000000010000100100000010101010010000001010101001000010010000000100001000000000000000000000000000000000000000",
"00011111000111110001111100001111000011110000000000010100100100001010101010011111000111110001111100001111000000000000010000010100100000000001000010011111000100001001111100011111000000000000101000010000100100001000000000011111000111110010101010011111001010101001111100011111000111110000000000000000000000000000000000000000",
"00010000000100100001000000000000100000001000000000010010100100001010010010010000100100000001001000000000100000000000010000010010100000000001000010010010000100001001000000010010000000000000010000010000100100001000000000010010000100000010010010010000001001001001000010010000000100100000000000000000000000000000000000000000",
"00010000000100010001000000010000100100001000000000010010100100001010010010010000100100000001000100010000100000000000010000010010100000000001000010010001000100001001000000010001000000000000010000010000100100001000000000010001000100000010010010010000001001001001000010010000000100010000000000000000000000000000000000000000",
"00010000000100001001111110001111000011110000000000010000100011110010000010011111000111111001000010001111000000000001111100010000100000000000111100010000100111100001111110010000100000000000010000001111000011110000000000010000100111111010000010011111101000001001111100011111100100001000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
"00000011110000010000010000011110000000011110000001111100001111111000000111100001111110001111111100111111100111100000000000001100011100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00001100001000010000010001100001100001100001100010000010001000000000001000010001000001001000000000100000000100010000000000010100100010010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00010000000100010000010010000000010010000000010010000000001000000000001000000001000001001000000000100000000100001000000000100100100010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00010000000000010000010010000000010010000000010001111100001111100000000111110001000001001111110000111110000100001000000000000100000100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00010000000000011111110010000000010010000000010000000010001000000000000000001001111110001000000000100000000100001001110000000100001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00010000000100010000010010000000010010000000010010000010001000000000001000001001000000001000000000100000000100001000000000000100010000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00001100001000010000010001100001100001100001100001000010001000000000000100001001000000001000000000100000000100010000000000000100111110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000011110000010000010000011110000000011110000000111100001111111000000011110001000000001111111100111111100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'),
(others => '0'));

signal rom_numbers: pamet_nmb := (
"00000000000000000000000000000000",
"00000001111111111111110000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001000000000000010000000000",
"00000001111111111111110000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000001110000000000000",
"00000000000000011110000000000000",
"00000000000000111110000000000000",
"00000000000001101110000000000000",
"00000000000011001110000000000000",
"00000000000110001110000000000000",
"00000000000000001110000000000000",
"00000000000000001110000000000000",
"00000000000000001110000000000000",
"00000000000000001110000000000000",
"00000000000000001110000000000000",
"00000000000000001110000000000000",
"00000000000000001110000000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000001111110000000000000000",
"00000000110000001100000000000000",
"00000011000000000011000000000000",
"00000011000000000011000000000000",
"00000011000000000011000000000000",
"00000000000000001100000000000000",
"00000000000000110000000000000000",
"00000000000011000000000000000000",
"00000000001100000000000000000000",
"00000000110000000000000000000000",
"00000011000000000000000000000000",
"00000011111111111111000000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000001111111111110000000000",
"00000000110000000000001100000000",
"00000011000000000000000011000000",
"00000011000000000000000011000000",
"00000000000000000000000011000000",
"00000000000000000000000011000000",
"00000000000011111111111100000000",
"00000000000000000000000011000000",
"00000000000000000000000011000000",
"00000011000000000000000011000000",
"00000011000000000000000011000000",
"00000000110000000000001100000000",
"00000000001111111111110000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000000000000011000000000000",
"00000000000000001100000000000000",
"00000000000000110000000000000000",
"00000000000011000000000000000000",
"00000000001100000000110000000000",
"00000000110000000000110000000000",
"00000011000000000000110000000000",
"00001111111111111111111111110000",
"00000000000000000000110000000000",
"00000000000000000000110000000000",
"00000000000000000000110000000000",
"00000000000000000000110000000000",
"00000000000000000000110000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000001111111111111111000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001111111111111111000000000",
"00000000000000000000001000000000",
"00000000000000000000001000000000",
"00000000000000000000001000000000",
"00000000000000000000001000000000",
"00000011111111111111111000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000001111111111111111111000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001000000000000000000000000",
"00000001111111111111111111000000",
"00000001000000000000000001000000",
"00000001000000000000000001000000",
"00000001000000000000000001000000",
"00000001000000000000000001000000",
"00000001111111111111111111000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000011111111111111110000000",
"00000000000000000000001110000000",
"00000000000000000000011000000000",
"00000000000000000000110000000000",
"00000000000000000011100000000000",
"00000000000111111111111100000000",
"00000000000000011100000000000000",
"00000000000000110000000000000000",
"00000000000001100000000000000000",
"00000000000111000000000000000000",
"00000000001100000000000000000000",
"00000000011000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000000011111111100000000000",
"00000000001100000000011000000000",
"00000000001000000000001000000000",
"00000000001000000000001000000000",
"00000000001000000000001000000000",
"00000000000111111111110000000000",
"00000000000110000000110000000000",
"00000000011000000000001100000000",
"00000000010000000000000100000000",
"00000000010000000000000100000000",
"00000000010000000000000100000000",
"00000000001100000000011000000000",
"00000000000011111111100000000000",
"00000000000000000000000000000000",
(others => '0'),
"00000000000000000000000000000000",
"00000000111111111111111100000000",
"00000000100000000000000100000000",
"00000000100000000000000100000000",
"00000000100000000000000100000000",
"00000000100000000000000100000000",
"00000000111111111111111100000000",
"00000000000000000000000100000000",
"00000000000000000000000100000000",
"00000000000000000000000100000000",
"00000000000000000000000100000000",
"00000000000000000000000100000000",
"00000000000000000000000100000000",
"00000000000000000000000100000000",
"00000000000000000000000000000000",
     (others => '0')
	  );
  
	signal sx : std_logic_vector(11 downto 0) := "000001000000";
	signal diffx : std_logic_vector(11 downto 0);
  
  
	--KEYBOARD
	signal kbrd_data_out : std_logic_vector(15 downto 0);
	signal kbrd_data_vld : std_logic;
	signal kbrd_data_vld_last : std_logic := '1';
	--signal kbrd_waiting : std_logic := '1';
	--signal kbrd_waiter : integer range 0 to 100001;

	signal pressed_button_index: integer range 0 to 17 := 17; -- 17 == nezm��knut� nic
	signal dir_lr : std_logic := '1';

	signal cntbg1 : std_logic_vector(3 downto 0);
	signal cntbg2 : std_logic_vector(3 downto 0);
	signal cntbg3 : std_logic_vector(3 downto 0);

begin

-- entity �asova��
gen_1mhz: entity work.engen generic map ( MAXVALUE => 39) port map ( CLK => CLK, ENABLE => '1', EN => en_1MHz );
gen_20hz: entity work.engen generic map ( MAXVALUE => 12500) port map ( CLK => CLK, ENABLE => en_1MHz, EN => en_20Hz );
--gen_1hz: entity work.engen generic map ( MAXVALUE => 10) port map ( CLK => CLK, ENABLE => en_20Hz, EN => en_1Hz );
gen_2hz: entity work.engen generic map ( MAXVALUE => 20) port map ( CLK => CLK, ENABLE => en_20Hz, EN => en_2Hz );
gen_4hz: entity work.engen generic map ( MAXVALUE => 40) port map ( CLK => CLK, ENABLE => en_20Hz, EN => en_4Hz );
gen_8hz: entity work.engen generic map ( MAXVALUE => 80) port map ( CLK => CLK, ENABLE => en_20Hz, EN => en_8Hz );
gen_16hz: entity work.engen generic map ( MAXVALUE => 160) port map ( CLK => CLK, ENABLE => en_20Hz, EN => en_16Hz );

-- entita pro generov�n� random ��sel, viz je�t� defaultn� nastaven� random_nmb
random_1: entity work.random port map( CLK => clk, RANDOM_NMB => random_nmb );

-- entita VGA
vga: entity work.vga_controller(arch_vga_controller)
  port map(
    CLK => CLK,
    RST => RESET,
    ENABLE => '1',
    MODE => vga_mode,
    DATA_RED => red,
    DATA_GREEN => green,
    DATA_BLUE => blue,
    ADDR_COLUMN => vgaCol,
    ADDR_ROW => vgaRow,
    VGA_RED => RED_V,
    VGA_GREEN => GREEN_V,
    VGA_BLUE => BLUE_V,
    VGA_HSYNC => HSYNC_V,
    VGA_VSYNC => VSYNC_V
  );

-- entita kl�vesnice  
	kbrd_ctrl: entity work.keyboard_controller(arch_keyboard)
	generic map (READ_INTERVAL => 1000000)
	port map (
		CLK => CLK,
		RST => RESET,

		DATA_OUT => kbrd_data_out(15 downto 0),
		DATA_VLD => kbrd_data_vld,
   
		KB_KIN   => KIN,
		KB_KOUT  => KOUT
	);
	
-- nastaven� m�du obrazovky  
setmode(r640x480x60, vga_mode);

process (CLK,random_nmb)
	variable temp : integer := 0;
	variable max_current_nmb_index : integer := 1;
begin
	if ( CLK'event ) and ( CLK = '1' ) then
		temp := conv_integer(random_nmb(2 downto 0))+conv_integer(random_nmb(3))+conv_integer(random_nmb(4))+conv_integer(random_nmb(5));
	
		if(kbrd_data_vld = '1') then
			key_pressed <= NONE;
				case kbrd_data_out is
					when "0000000000000001" => key_pressed <= K1; 		number_pressed <= "0001";
					when "0000000000000010" => key_pressed <= K4; 		number_pressed <= "0100";
					when "0000000000000100" => key_pressed <= K7; 		number_pressed <= "0111";
					when "0000000000001000" => key_pressed <= KSTAR; 	number_pressed <= "1111";
					when "0000000000010000" => key_pressed <= K2;		number_pressed <= "0010";
					when "0000000000100000" => key_pressed <= K5;		number_pressed <= "0101";
					when "0000000001000000" => key_pressed <= K8;		number_pressed <= "1000";
					when "0000000010000000" => key_pressed <= K0;		number_pressed <= "0000";
					when "0000000100000000" => key_pressed <= K3;		number_pressed <= "0011";
					when "0000001000000000" => key_pressed <= K6;		number_pressed <= "0110";
					when "0000010000000000" => key_pressed <= K9;		number_pressed <= "1001";
					when "0000100000000000" => key_pressed <= KHASH; 	number_pressed <= "1111";
					when "0001000000000000" => key_pressed <= KA; 		number_pressed <= "1111";
					when "0010000000000000" => key_pressed <= KB; 		number_pressed <= "1111";
					when "0100000000000000" => key_pressed <= KC;		number_pressed <= "1111";
					when "1000000000000000" => key_pressed <= KD;		number_pressed <= "1111";
					when others => key_pressed <= NONE;
				end case;
		else
			key_pressed <= NONE;
		end if;

		case game_state is
			-- generace ��sel
			when WELCOME_SCREEN =>
				if(key_pressed = KHASH ) then
					current_nmb_index <= MIN_INDEX;
					game_state <= GEN_NMB;
				elsif(key_pressed = KA)then
					game_state <= CONFIG_SPEED;
				end if;
			when CONFIG_SPEED =>
				-- konfigurace rychlosti zobrazov�n� n�hodn�ch ��slic
				if(key_pressed = K1 ) then
					game_speed <= "100";
					game_state <= CONFIG_SPEED;
				elsif(key_pressed = K2)then
					game_speed <= "010";
					game_state <= CONFIG_SPEED;
				elsif(key_pressed = K3)then
					game_speed <= "001";
					game_state <= CONFIG_SPEED;
				elsif(key_pressed = KSTAR)then
					game_state <= WELCOME_SCREEN;
				end if;
			when WAITING_SCREEN =>
				current_nmb_index <= MIN_INDEX;
				game_state <= GEN_NMB;
			when GEN_NMB =>
				--if (current_nmb_index = temp) then
				--	generated_rand(current_nmb_index) <= 1;
				--else
				generated_rand(current_nmb_index) <= temp;
				-- nastaven� neopakov�n�!!!
				--	end if;
				if(current_nmb_index = MAX_INDEX) then
					game_state <= SHOWING_NUMBERS;
					current_nmb_index <= MIN_INDEX;
				else 
					current_nmb_index <= current_nmb_index+1;
				end if;
			when SHOWING_NUMBERS =>
				-- game - zobrazuje ��sla pro zapamatov�n�
				if( (en_4Hz = '1' and game_speed(0) = '1') or (en_8Hz = '1' and game_speed(1) = '1') or (en_16Hz = '1' and game_speed(2) = '1')) then
					if(current_nmb_index /= MAX_INDEX) then
						current_nmb_index <= current_nmb_index + 1;
					end if;
				end if; 
				max_current_nmb_index := game_level+2;
				if( current_nmb_index = MAX_INDEX OR current_nmb_index >= max_current_nmb_index) then -- OR current_nmb_index > conv_integer(game_level)
					current_nmb_index <= MIN_INDEX;
					text <= BEFORE_WRITING_NUMBERS;
					number_pressed <= "1111";
					game_state <= WRITING_NUMBERS;
				end if;

			when WRITING_NUMBERS =>
					-- playing - zad�v�n� ��sel
					if( en_4Hz = '1' ) then
						if ( key_pressed = KD) then
							game_state <= LEVEL_END_OK;
						end if;
						max_current_nmb_index := game_level+2;
						if ( current_nmb_index >= max_current_nmb_index ) then
							-- level acomplished
							game_state <= LEVEL_END_OK;
							text <= LEVEL_OK;
							if(game_level = MAX_INDEX) then 
								game_level <= 1;
							else
								game_level <= game_level+1;
							end if;
							max_current_nmb_index := game_level+2;
							current_nmb_index <= MIN_INDEX;
						elsif (key_pressed = KA) then
							game_state <= SHOWING_NUMBERS;
							current_nmb_index <= MIN_INDEX;
						else 
								if(conv_integer(number_pressed) /= conv_integer(generated_rand(current_nmb_index)) and number_pressed /= "1111") then
										-- nesouhlas� vysko�� z levelu na 
										number_pressed <= "1111";
										game_state <= LEVEL_END_BAD;
										text <= LEVEL_BAD;
								elsif ( number_pressed /= "1111") then
									if ( current_nmb_index = MAX_INDEX ) then
										current_nmb_index <= MIN_INDEX;
									else
										current_nmb_index <= current_nmb_index +1;
									end if;
									number_pressed <= "1111";
								end if;
						end if;
					end if;
				--end if;
			when LEVEL_END_BAD =>
				if (text = LEVEL_BAD) then
					if(key_pressed = KSTAR) then
						-- p�ejde na start - nastav�m defaultn� hodnoty a p�enastav�m game_state na init
						game_state <= WELCOME_SCREEN;
						text <= NONE;
					end if;
				end if;
				-- �sp�n� ukon�en� levelu
			when LEVEL_END_OK =>
				if(key_pressed = KSTAR) then
					current_nmb_index <= MIN_INDEX;
					game_state <= GEN_NMB;
				end if;
				
				--if (text = LEVEL_OK) then
					--if(key_pressed = KHASH) then
						-- p�ejde na dal�� level - zv���m level value a game_state na generov�n� ��sel
						--game_state <= GEN_NMB;
						--text <= NONE;
					--end if;
				--end if;
				-- ne�sp�n� ukon�en� levelu
		end case;
   end if;
end process;

-- type t_game_states is (INIT,WELCOME_SCREEN,WAITING_SCREEN,GEN_NMB, SHOWING_NUMBERS, WRITING_NUMBERS,WAITING_FOR_KEY,LEVEL_END_BAD,LEVEL_END_OK);

rgb <= "111"&"111"&"111" when game_state = SHOWING_NUMBERS and rom_numbers(16*generated_rand(current_nmb_index)+conv_integer(vgaRow(3 downto 0)) )(conv_integer(vgaCol(4 downto 0)))='1' else 
		 "111"&"111"&"111" when game_state = WRITING_NUMBERS and number_pressed /= "1111" and rom_numbers(16*conv_integer(number_pressed)+conv_integer(vgaRow(3 downto 0)))(conv_integer(vgaCol(4 downto 0)))='1' else 
		 "000"&"000"&"000";

rgbMsg <= "111"&"111"&"111" when ( game_state = WELCOME_SCREEN OR game_state = GEN_NMB ) and rom_msg(conv_integer(vgaRow(2 downto 0)))(conv_integer(vgaCol(8 downto 0))-100)='1' else 
			 "000"&"111"&"000" when game_state = LEVEL_END_OK and rom_msg(16*1 + conv_integer(vgaRow(2 downto 0)))(conv_integer(vgaCol(8 downto 0))-100)='1' else 
			 "111"&"000"&"000" when game_state = LEVEL_END_BAD and rom_msg(16*2 + conv_integer(vgaRow(2 downto 0)))(conv_integer(vgaCol(8 downto 0))-100)='1' else 
			 "111"&"111"&"111" when game_state = WRITING_NUMBERS and rom_msg(16*3 + conv_integer(vgaRow(2 downto 0)))(conv_integer(vgaCol(8 downto 0))-100)='1' else 
			 "111"&"111"&"111" when game_state = CONFIG_SPEED and rom_msg(16*4 + conv_integer(vgaRow(2 downto 0)))(conv_integer(vgaCol(8 downto 0))-100)='1' else 
			 "000"&"000"&"000";

rgbLvlMsg <= "111"&"111"&"111" when ( game_state /= WELCOME_SCREEN) and rom_lvl(conv_integer(vgaRow(2 downto 0)))(conv_integer(vgaCol(4 downto 0)))='1' else 
      "000"&"000"&"000";
		 
rgbLvlNmb <= "111"&"111"&"111" when ( game_state /= WELCOME_SCREEN) and rom_numbers(game_level*16+conv_integer(vgaRow(3 downto 0)))(conv_integer(vgaCol(4 downto 0)))='1' else 
       "000"&"000"&"000";
		 
rgbf <= 	
			rgb 			when (vgaRow(11 downto 4) = "00010000") and (vgaCol(11 downto 5) = "0001000")  else
			"000"&"111"&"000" when game_speed(0) = '1' and game_state = CONFIG_SPEED and (vgaRow(11 downto 0) = "000000101111") and vgaCol(11 downto 2) = "00111011" else --and vgaCol(7 downto 3) = "1111" else
			"000"&"111"&"000" when game_speed(1) = '1' and game_state = CONFIG_SPEED and (vgaRow(11 downto 0) = "000000101111") and vgaCol(11 downto 2) = "00111001" else -- and vgaCol(7 downto 3) = "1011" else
			"000"&"111"&"000" when game_speed(2) = '1' and game_state = CONFIG_SPEED and (vgaRow(11 downto 0) = "000000101111") and vgaCol(11 downto 2) = "00111000" else --and vgaCol(7 downto 3) = "1001" else
			rgbMsg 		when (vgaRow(11 downto 3) = "000000101") and conv_integer(vgaCol) > 100 and conv_integer(vgaCol) < 500 else --and (vgaCol(11 downto 7) = "00000")
			rgbLvlMsg	when (vgaRow(11 downto 3) = "000001111") and conv_integer(vgaCol) > 194 and conv_integer(vgaCol) < 235 else
			rgbLvlNmb	when (vgaRow(11 downto 4) = "00000111") and conv_integer(vgaCol) > 255 and conv_integer(vgaCol) < 285 else
			"000"&"000"&"000";

red <= rgbf(8 downto 6);
green <= rgbf(5 downto 3);
blue <= rgbf(2 downto 0);
end;